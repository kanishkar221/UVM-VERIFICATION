UVM_INFO env.sv(10) @ 0: uvm_test_top.env [ENV] Environment Created
UVM_INFO sequence.sv(11) @ 0: uvm_test_top.env.agent.sequencer@@seq [SEQ] Sequence Starts
UVM_INFO scoreboard.sv(29) @ 6: uvm_test_top.env.sb [SB] PASS ---> Input:clk=0  wr=0  d_in=0  addr=0  Actual Output: d_out=0 || Expected Output: exp_d_out=0
UVM_INFO scoreboard.sv(23) @ 16: uvm_test_top.env.sb [SB] WRITE PASS -----> Input:clk=0  wr=1  d_in=155 addr=9  d_out=0
UVM_INFO scoreboard.sv(23) @ 26: uvm_test_top.env.sb [SB] WRITE PASS -----> Input:clk=0  wr=1  d_in=0 addr=3  d_out=0
UVM_INFO scoreboard.sv(29) @ 36: uvm_test_top.env.sb [SB] PASS ---> Input:clk=0  wr=0  d_in=11  addr=4  Actual Output: d_out=0 || Expected Output: exp_d_out=0
UVM_INFO scoreboard.sv(23) @ 46: uvm_test_top.env.sb [SB] WRITE PASS -----> Input:clk=0  wr=1  d_in=188 addr=5  d_out=0
UVM_INFO scoreboard.sv(23) @ 56: uvm_test_top.env.sb [SB] WRITE PASS -----> Input:clk=0  wr=1  d_in=251 addr=4  d_out=0
UVM_INFO scoreboard.sv(29) @ 66: uvm_test_top.env.sb [SB] PASS ---> Input:clk=0  wr=0  d_in=200  addr=2  Actual Output: d_out=0 || Expected Output: exp_d_out=0
UVM_INFO scoreboard.sv(23) @ 76: uvm_test_top.env.sb [SB] WRITE PASS -----> Input:clk=0  wr=1  d_in=58 addr=6  d_out=0
UVM_INFO scoreboard.sv(23) @ 86: uvm_test_top.env.sb [SB] WRITE PASS -----> Input:clk=0  wr=1  d_in=221 addr=2  d_out=0
UVM_INFO scoreboard.sv(23) @ 96: uvm_test_top.env.sb [SB] WRITE PASS -----> Input:clk=0  wr=1  d_in=14 addr=8  d_out=0
UVM_INFO scoreboard.sv(29) @ 106: uvm_test_top.env.sb [SB] PASS ---> Input:clk=0  wr=0  d_in=229  addr=9  Actual Output: d_out=155 || Expected Output: exp_d_out=155
UVM_INFO scoreboard.sv(23) @ 116: uvm_test_top.env.sb [SB] WRITE PASS -----> Input:clk=0  wr=1  d_in=74 addr=8  d_out=155
UVM_INFO scoreboard.sv(29) @ 126: uvm_test_top.env.sb [SB] PASS ---> Input:clk=0  wr=0  d_in=223  addr=7  Actual Output: d_out=0 || Expected Output: exp_d_out=0
UVM_INFO scoreboard.sv(29) @ 136: uvm_test_top.env.sb [SB] PASS ---> Input:clk=0  wr=0  d_in=120  addr=4  Actual Output: d_out=251 || Expected Output: exp_d_out=251
UVM_INFO scoreboard.sv(29) @ 146: uvm_test_top.env.sb [SB] PASS ---> Input:clk=0  wr=0  d_in=88  addr=2  Actual Output: d_out=221 || Expected Output: exp_d_out=221
UVM_INFO scoreboard.sv(23) @ 156: uvm_test_top.env.sb [SB] WRITE PASS -----> Input:clk=0  wr=1  d_in=175 addr=4  d_out=221
UVM_INFO scoreboard.sv(29) @ 166: uvm_test_top.env.sb [SB] PASS ---> Input:clk=0  wr=0  d_in=78  addr=10  Actual Output: d_out=0 || Expected Output: exp_d_out=0
UVM_INFO scoreboard.sv(23) @ 176: uvm_test_top.env.sb [SB] WRITE PASS -----> Input:clk=0  wr=1  d_in=240 addr=0  d_out=0
UVM_INFO scoreboard.sv(29) @ 186: uvm_test_top.env.sb [SB] PASS ---> Input:clk=0  wr=0  d_in=195  addr=5  Actual Output: d_out=188 || Expected Output: exp_d_out=188
UVM_INFO scoreboard.sv(29) @ 196: uvm_test_top.env.sb [SB] PASS ---> Input:clk=0  wr=0  d_in=130  addr=2  Actual Output: d_out=221 || Expected Output: exp_d_out=221
