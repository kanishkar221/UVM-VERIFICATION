interface FA_if;
  logic a;
  logic b;
  logic cin;
  logic sum;
  logic cout;
endinterface  
