UVM_INFO env.sv(10) @ 0: uvm_test_top.env [ENV] Environment Created
UVM_INFO sequence.sv(11) @ 0: uvm_test_top.env.agent.sequencer@@seq [SEQ] Sequence Starts
UVM_INFO scoreboard.sv(29) @ 6: uvm_test_top.env.sb [SB] PASS ---> Input:clk=0  wr=0  d_in=0  addr=0  Actual Output: d_out=0 || Expected Output: exp_d_out=0
UVM_INFO scoreboard.sv(23) @ 16: uvm_test_top.env.sb [SB] WRITE PASS -----> Input:clk=0  wr=1  d_in=155 addr=9  d_out=0
UVM_INFO scoreboard.sv(23) @ 26: uvm_test_top.env.sb [SB] WRITE PASS -----> Input:clk=0  wr=1  d_in=0 addr=3  d_out=0
UVM_INFO scoreboard.sv(29) @ 36: uvm_test_top.env.sb [SB] PASS ---> Input:clk=0  wr=0  d_in=11  addr=4  Actual Output: d_out=0 || Expected Output: exp_d_out=0
UVM_INFO scoreboard.sv(23) @ 46: uvm_test_top.env.sb [SB] WRITE PASS -----> Input:clk=0  wr=1  d_in=188 addr=5  d_out=0
UVM_INFO scoreboard.sv(23) @ 56: uvm_test_top.env.sb [SB] WRITE PASS -----> Input:clk=0  wr=1  d_in=251 addr=4  d_out=0
UVM_INFO scoreboard.sv(29) @ 66: uvm_test_top.env.sb [SB] PASS ---> Input:clk=0  wr=0  d_in=200  addr=2  Actual Output: d_out=0 || Expected Output: exp_d_out=0
UVM_INFO scoreboard.sv(23) @ 76: uvm_test_top.env.sb [SB] WRITE PASS -----> Input:clk=0  wr=1  d_in=58 addr=6  d_out=0
UVM_INFO scoreboard.sv(23) @ 86: uvm_test_top.env.sb [SB] WRITE PASS -----> Input:clk=0  wr=1  d_in=221 addr=2  d_out=0
UVM_INFO scoreboard.sv(23) @ 96: uvm_test_top.env.sb [SB] WRITE PASS -----> Input:clk=0  wr=1  d_in=14 addr=8  d_out=0
