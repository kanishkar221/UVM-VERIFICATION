interface counter_if;
  logic clk;
  logic reset;
  logic enable;
  logic [3:0] count;
endinterface
  
