UVM_INFO env.sv(10) @ 0: uvm_test_top.env [ENV] Environment Created
UVM_INFO sequence.sv(11) @ 0: uvm_test_top.env.agent.sequencer@@seq [SEQ] Sequence starts
UVM_INFO scoreboard.sv(29) @ 6: uvm_test_top.env.sb [SB] PASS ----> reset=1  enable=0  Actual count=0  Expected count=0
----------------------------------------------------------------
UVM_INFO scoreboard.sv(29) @ 16: uvm_test_top.env.sb [SB] PASS ----> reset=0  enable=1  Actual count=1  Expected count=1
----------------------------------------------------------------
UVM_INFO scoreboard.sv(29) @ 26: uvm_test_top.env.sb [SB] PASS ----> reset=0  enable=0  Actual count=1  Expected count=1
----------------------------------------------------------------
UVM_INFO scoreboard.sv(29) @ 36: uvm_test_top.env.sb [SB] PASS ----> reset=0  enable=1  Actual count=2  Expected count=2
----------------------------------------------------------------
UVM_INFO scoreboard.sv(29) @ 46: uvm_test_top.env.sb [SB] PASS ----> reset=0  enable=0  Actual count=2  Expected count=2
----------------------------------------------------------------
UVM_INFO scoreboard.sv(29) @ 56: uvm_test_top.env.sb [SB] PASS ----> reset=0  enable=0  Actual count=2  Expected count=2
----------------------------------------------------------------
UVM_INFO scoreboard.sv(29) @ 66: uvm_test_top.env.sb [SB] PASS ----> reset=0  enable=0  Actual count=2  Expected count=2
----------------------------------------------------------------
UVM_INFO scoreboard.sv(29) @ 76: uvm_test_top.env.sb [SB] PASS ----> reset=0  enable=0  Actual count=2  Expected count=2
----------------------------------------------------------------
UVM_INFO scoreboard.sv(29) @ 86: uvm_test_top.env.sb [SB] PASS ----> reset=0  enable=0  Actual count=2  Expected count=2
----------------------------------------------------------------
UVM_INFO scoreboard.sv(29) @ 96: uvm_test_top.env.sb [SB] PASS ----> reset=0  enable=1  Actual count=3  Expected count=3
----------------------------------------------------------------
UVM_INFO scoreboard.sv(29) @ 106: uvm_test_top.env.sb [SB] PASS ----> reset=0  enable=1  Actual count=4  Expected count=4
----------------------------------------------------------------
UVM_INFO scoreboard.sv(29) @ 116: uvm_test_top.env.sb [SB] PASS ----> reset=0  enable=1  Actual count=5  Expected count=5
----------------------------------------------------------------
UVM_INFO scoreboard.sv(29) @ 126: uvm_test_top.env.sb [SB] PASS ----> reset=0  enable=1  Actual count=6  Expected count=6
----------------------------------------------------------------
UVM_INFO scoreboard.sv(29) @ 136: uvm_test_top.env.sb [SB] PASS ----> reset=0  enable=1  Actual count=7  Expected count=7
----------------------------------------------------------------
UVM_INFO scoreboard.sv(29) @ 146: uvm_test_top.env.sb [SB] PASS ----> reset=0  enable=1  Actual count=8  Expected count=8
----------------------------------------------------------------
UVM_INFO scoreboard.sv(29) @ 156: uvm_test_top.env.sb [SB] PASS ----> reset=0  enable=1  Actual count=9  Expected count=9
----------------------------------------------------------------
