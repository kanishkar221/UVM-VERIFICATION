UVM_INFO FA_env.sv(10) @ 0: uvm_test_top.env [ENV] Environment Created
UVM_INFO FA_sequence.sv(11) @ 0: uvm_test_top.env.agent.sequencer@@seq [SEQ] Sequence starts
UVM_INFO FA_scoreboard.sv(25) @ 10: uvm_test_top.env.sb [SB] PASS----> INPUT:a=0 | b=0 | cin=1 | Actual output: sum=1 | cout=0 || Expected output:sum=1 |cout=0
UVM_INFO FA_scoreboard.sv(25) @ 20: uvm_test_top.env.sb [SB] PASS----> INPUT:a=0 | b=0 | cin=1 | Actual output: sum=1 | cout=0 || Expected output:sum=1 |cout=0
UVM_INFO FA_scoreboard.sv(25) @ 30: uvm_test_top.env.sb [SB] PASS----> INPUT:a=0 | b=1 | cin=1 | Actual output: sum=0 | cout=1 || Expected output:sum=0 |cout=1
UVM_INFO FA_scoreboard.sv(25) @ 40: uvm_test_top.env.sb [SB] PASS----> INPUT:a=1 | b=0 | cin=1 | Actual output: sum=0 | cout=1 || Expected output:sum=0 |cout=1
UVM_INFO FA_scoreboard.sv(25) @ 50: uvm_test_top.env.sb [SB] PASS----> INPUT:a=1 | b=1 | cin=1 | Actual output: sum=1 | cout=1 || Expected output:sum=1 |cout=1
UVM_INFO FA_scoreboard.sv(25) @ 60: uvm_test_top.env.sb [SB] PASS----> INPUT:a=0 | b=0 | cin=1 | Actual output: sum=1 | cout=0 || Expected output:sum=1 |cout=0
UVM_INFO FA_scoreboard.sv(25) @ 70: uvm_test_top.env.sb [SB] PASS----> INPUT:a=1 | b=1 | cin=1 | Actual output: sum=1 | cout=1 || Expected output:sum=1 |cout=1
UVM_INFO FA_scoreboard.sv(25) @ 80: uvm_test_top.env.sb [SB] PASS----> INPUT:a=0 | b=0 | cin=0 | Actual output: sum=0 | cout=0 || Expected output:sum=0 |cout=0
UVM_INFO FA_scoreboard.sv(25) @ 90: uvm_test_top.env.sb [SB] PASS----> INPUT:a=1 | b=0 | cin=1 | Actual output: sum=0 | cout=1 || Expected output:sum=0 |cout=1
