UVM_INFO ha_env.sv(10) @ 0: uvm_test_top.env [ENV] Environment Created
UVM_INFO ha_sequence.sv(11) @ 0: uvm_test_top.env.agent.sequencer@@seq [SEQ] Sequence starts
UVM_INFO ha_scoreboard.sv(24) @ 10: uvm_test_top.env.sb [SB] PASS----> INPUT:a=0 | b=0 | Actual output: sum=0 | carry=0 || Expected output:sum=0 | carry=0
UVM_INFO ha_scoreboard.sv(24) @ 20: uvm_test_top.env.sb [SB] PASS----> INPUT:a=0 | b=1 | Actual output: sum=1 | carry=0 || Expected output:sum=1 | carry=0
UVM_INFO ha_scoreboard.sv(24) @ 30: uvm_test_top.env.sb [SB] PASS----> INPUT:a=0 | b=1 | Actual output: sum=1 | carry=0 || Expected output:sum=1 | carry=0
UVM_INFO ha_scoreboard.sv(24) @ 40: uvm_test_top.env.sb [SB] PASS----> INPUT:a=1 | b=1 | Actual output: sum=0 | carry=1 || Expected output:sum=0 | carry=1
UVM_INFO ha_scoreboard.sv(24) @ 50: uvm_test_top.env.sb [SB] PASS----> INPUT:a=1 | b=0 | Actual output: sum=1 | carry=0 || Expected output:sum=1 | carry=0
UVM_INFO ha_scoreboard.sv(24) @ 60: uvm_test_top.env.sb [SB] PASS----> INPUT:a=0 | b=1 | Actual output: sum=1 | carry=0 || Expected output:sum=1 | carry=0
UVM_INFO ha_scoreboard.sv(24) @ 70: uvm_test_top.env.sb [SB] PASS----> INPUT:a=1 | b=0 | Actual output: sum=1 | carry=0 || Expected output:sum=1 | carry=0
UVM_INFO ha_scoreboard.sv(24) @ 80: uvm_test_top.env.sb [SB] PASS----> INPUT:a=0 | b=1 | Actual output: sum=1 | carry=0 || Expected output:sum=1 | carry=0
UVM_INFO ha_scoreboard.sv(24) @ 90: uvm_test_top.env.sb [SB] PASS----> INPUT:a=1 | b=0 | Actual output: sum=1 | carry=0 || Expected output:sum=1 | carry=0
